entity eighteenBitRow is 
	
	port (
	
	);
	
end eighteenBitRow;

architecture rtl of eighteenBitRow is 

	component oneBitAdder 
		port (		
		i_CarryIn		: IN	STD_LOGIC;
		i_Ai, i_Bi		: IN	STD_LOGIC;
		o_Sum, o_CarryOut	: OUT	STD_LOGIC);

	begin 
	
	
	
	
end rtl; 